module registerFile (
    input logic [9:0] D,
    input logic ENW, ENRO, ENR1, CLKb,
    input logic [2:0] WRA, RDA0, RDA1,
    output logic [9:0] Q0, Q1
);




endmodule