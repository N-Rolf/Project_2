//top level file for 10-bit processor
module ARM_processor (
    input logic 
    output logic
);



endmodule