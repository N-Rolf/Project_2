module ARM_processor (
    input logic 
    output logic
);



endmodule